module top_module( output one );

// Insert your code here
    assign one = 'b1;

endmodule
